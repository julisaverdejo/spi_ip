module spi_ip(
);

endmodule